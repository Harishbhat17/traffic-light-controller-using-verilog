`timescale 1ns / 1ps
module pro1(output reg [3:0] red,yel,gre,input clk,rst);
parameter s0=3'b000,s1=3'b001,s2=3'b010,s3=3'b011,s4=3'b100;
reg [2:0]ns,cs;
reg [5:0] counter;

always @(posedge clk,posedge rst)
begin
if(rst)
begin
cs<=s0;
counter<=0;
end
else
begin
cs<=ns;
counter<=counter+6'b000001;
end
end
always@(*)
begin
case(cs)
s0:
ns<=s1; 
s1:
if(counter >=16)
begin
ns<=s2; 
end
else
ns<=s1;
s2:
if(counter >=24)
begin
ns<=s3; 
end 
else
ns<=s2;
s3:
if(counter >=32)
begin
ns<=s4; 
end 
else
ns<=s3;
s4:
if(counter>=40)begin
counter<=0;
ns=s1;
end 
else
ns=s1;
endcase
end
always@(ns,cs)
begin
case(cs)
s0:
begin
red<=4'b0000;
yel<=4'b0000;
gre<=4'b0000;
end 
s1:
if(counter<12)
begin
red<=4'b1010;
yel<=4'b0000;
gre<=4'b0101;
end 
else
begin
red<=4'b0000;
yel<=4'b0101;
gre<=4'b1010;
end
s2:
if(counter<18)
begin
red<=4'b0101;
yel<=4'b0000;
gre<=4'b1010;
end 
else
begin
red<=4'b0000;
yel<=4'b0101;
gre<=4'b1010;
end
s3:
if(counter<24)
begin
red<=4'b1010;
yel<=4'b0000;
gre<=4'b0101;
end 
else
begin
red<=4'b0000;
yel<=4'b0101;
gre<=4'b1010;
end
s4:
if(counter<30)
begin
red<=4'b0101;
yel<=4'b0000;
gre<=4'b1010;
end 
else
begin
red<=4'b0000;
yel<=4'b0101;
gre<=4'b1010;
end
endcase
end
endmodule
